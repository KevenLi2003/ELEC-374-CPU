`timescale 1ns/10ps
module and_tb;

    // Control signals
    reg PCout, Zlowout, MDRout, R3out, R7out;
    reg MARin, Zin, PCin, MDRin, IRin, Yin;
    reg IncPC, Read, R3in, R4in, R7in;
    reg Clock;
    reg [31:0] Mdatain;

    // ALU control signal for AND operation
    reg [3:0] ALU_control;

    // States for FSM
    parameter Default = 4'b0000, Reg_load1a = 4'b0001, Reg_load1b = 4'b0010, Reg_load2a = 4'b0011,
              Reg_load2b = 4'b0100, Reg_load3a = 4'b0101, Reg_load3b = 4'b0110, T0 = 4'b0111,
              T1 = 4'b1000, T2 = 4'b1001, T3 = 4'b1010, T4 = 4'b1011, T5 = 4'b1100;

    reg [3:0] Present_state = Default;

    // Instantiate the datapath module
    datapath DUT (
        .clk(Clock), .reset(1'b0),
        .PCout(PCout), .Zlowout(Zlowout), .MDRout(MDRout), .R3out(R3out), .R7out(R7out),
        .MARin(MARin), .Zin(Zin), .PCin(PCin), .MDRin(MDRin), .IRin(IRin), .Yin(Yin),
        .IncPC(IncPC), .Read(Read), .AND(AND),
        .R3in(R3in), .R4in(R4in), .R7in(R7in),
        .Mdatain(Mdatain),
        .ALU_control(ALU_control) // Connect ALU control directly
    );

    // Clock generation
    initial begin
        Clock = 0;
        forever #10 Clock = ~Clock; // 20ns clock period
    end

    // FSM: Control sequence for the AND operation
    always @(posedge Clock) begin
        case (Present_state)
            Default: Present_state = Reg_load1a;
            Reg_load1a: Present_state = Reg_load1b;
            Reg_load1b: Present_state = Reg_load2a;
            Reg_load2a: Present_state = Reg_load2b;
            Reg_load2b: Present_state = Reg_load3a;
            Reg_load3a: Present_state = Reg_load3b;
            Reg_load3b: Present_state = T0;
            T0: Present_state = T1;
            T1: Present_state = T2;
            T2: Present_state = T3;
            T3: Present_state = T4;
            T4: Present_state = T5;
        endcase
    end

    // Apply control signals for each state
    always @(Present_state) begin
        case (Present_state)
            Default: begin
                // Initialize signals
                PCout <= 0; Zlowout <= 0; MDRout <= 0; R3out <= 0; R7out <= 0;
                MARin <= 0; Zin <= 0; PCin <= 0; MDRin <= 0; IRin <= 0; Yin <= 0;
                IncPC <= 0; Read <= 0; ALU_control <= 4'b0000;
                R3in <= 0; R4in <= 0; R7in <= 0; Mdatain <= 32'h00000000;
            end

            // Load data into R3
            Reg_load1a: begin
                Mdatain <= 32'h00000022; // Value for R3
                Read <= 1; MDRin <= 1;
            end
            Reg_load1b: begin
                Read <= 0; MDRin <= 0;
                MDRout <= 1; R3in <= 1;
                #15 MDRout <= 0; R3in <= 0;
            end

            // Load data into R7
            Reg_load2a: begin
                Mdatain <= 32'h00000024; // Value for R7
                Read <= 1; MDRin <= 1;
            end
            Reg_load2b: begin
                Read <= 0; MDRin <= 0;
                MDRout <= 1; R7in <= 1;
                #15 MDRout <= 0; R7in <= 0;
            end

            // Load data into R4 (this will hold the AND result later)
            Reg_load3a: begin
                Mdatain <= 32'h00000028; // Value for R4
                Read <= 1; MDRin <= 1;
            end
            Reg_load3b: begin
                Read <= 0; MDRin <= 0;
                MDRout <= 1; R4in <= 1;
                #15 MDRout <= 0; R4in <= 0;
            end

            // Perform AND operation
            T0: begin
                PCout <= 1; MARin <= 1; IncPC <= 1; Zin <= 1;
            end
            T1: begin
                PCout <= 0; MARin <= 0; IncPC <= 0; Zin <= 0;
                Zlowout <= 1; PCin <= 1; Read <= 1; MDRin <= 1;
                Mdatain <= 32'h2A2B8000; // Opcode for "AND R4, R3, R7"
            end
            T2: begin
                Read <= 0; MDRin <= 0;
                MDRout <= 1; IRin <= 1;
            end
            T3: begin
                MDRout <= 0; IRin <= 0;
                R3out <= 1; Yin <= 1;
            end
            T4: begin
                R3out <= 0; Yin <= 0;
                R7out <= 1; ALU_control <= 4'b0010; // Activate AND operation
                Zin <= 1;
            end
            T5: begin
                R7out <= 0; Zin <= 0;
                Zlowout <= 1; R4in <= 1;
                #15 Zlowout <= 0; R4in <= 0; // Store result into R4
            end
        endcase
    end

endmodule